module registers ();

endmodule