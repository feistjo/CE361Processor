module d_mem()

endmodule