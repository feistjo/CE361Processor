// do shit here idk man
// needs adders, mux, extender
`include "lib/sram.v"
`include "lib/syncram.v"

module pc_branch(pc_in, imm16, nPC_sel, pc_out);
   input [31:0] pc_in;
   input [15:0] imm16;
   input 	nPC_sel;
   output [31:0] pc_out;

   

   

    

   
endmodule // fuck_around
