// do shit here idk man


module pc_branch(A, imm16, nPC_sel, pc_out);
   input [31:0] A;
   input [15:0] imm16;
   input 	nPC_sel;
   output [31:0] pc_out;

   

    

   
endmodule // fuck_around
