// do shit here idk man


module fuck_around(A, B, out)
    input [31:0] A;
    input [31:0] B;
    output [31:0] out;

    // weeeeeeeee



endmodule